//WRITEME: takes multiple fifos and syncronizes/concats